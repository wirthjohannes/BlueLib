package BlueLib;

import BlueLibTests :: *;
export BlueLibTests :: *;

import BlueLibNetwork :: *;
export BlueLibNetwork :: *;

import BlueLibUtils :: *;
export BlueLibUtils :: *;

import PacketParser :: *;
export PacketParser :: *;

import PacketSender :: *;
export PacketSender :: *;

import BlueLibFIFO :: *;
export BlueLibFIFO :: *;

import BlueLibXilinxPrimitives :: *;
export BlueLibXilinxPrimitives :: *;

import TestHelpers :: *;
export TestHelpers :: *;

import Logging :: *;
export Logging :: *;

endpackage
